/***********************************************************************
 * A SystemVerilog top-level netlist to connect testbench to DUT
 **********************************************************************/

module top;
  //timeunit 1ns/1ns;

  // user-defined types are defined in instr_register_pkg.sv
  import instr_register_pkg::*;

  // clock variables
  logic clk;
  logic test_clk;

  // interconnecting signals
  // logic          load_en;
  // logic          reset_n;
  // opcode_t       opcode;
  // operand_t      operand_a, operand_b;
  // address_t      write_pointer, read_pointer;
  // instruction_t  instruction_word;
  tb_ifc laborator4(.clk(test_clk));
    // .load_en(load_en),
    // .reset_n(reset_n),
    // .opcode(opcode),
    // .operand_a(operand_a), 
    // .operand_b(operand_b),
    // .write_pointer(write_pointer),
    // .read_pointer(read_pointer),
    // .instruction_word(instruction_word)

  // instantiate testbench and connect ports
  instr_register_test test (.test_laborator_4(laborator4));

  // instantiate design and connect ports
  instr_register dut (
    .clk(clk),
    .load_en(laborator4.load_en),
    .reset_n(laborator4.reset_n),
    .operand_a(laborator4.operand_a),
    .operand_b(laborator4.operand_b),
    .opcode(laborator4.opcode),
    .write_pointer(laborator4.write_pointer),
    .read_pointer(laborator4.read_pointer),
    .instruction_word(laborator4.instruction_word)
   );

  // clock oscillators
  initial begin
    clk <= 0;
    forever #5  clk = ~clk;
  end

  initial begin
    test_clk <=0;
    // offset test_clk edges from clk to prevent races between
    // the testbench and the design
    #4 forever begin
      #2ns test_clk = 1'b1;
      #8ns test_clk = 1'b0;
    end
  end

endmodule: top
